library verilog;
use verilog.vl_types.all;
entity pipelined_computer_vlg_vec_tst is
end pipelined_computer_vlg_vec_tst;
